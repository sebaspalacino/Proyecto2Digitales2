`include "fifo.v"
`include "demux_id.v"
`include "mux_dst.v"
`include "demux_t.v"
module pcie_trans#(parameter BITNUMBER = 6,
			parameter LENGTH = 4)(
    input [BITNUMBER-1:0] data_in,
    input clk,
    input reset,
    input push,
    input pop_D0,
    input pop_D1,
    output wire [BITNUMBER-1:0] data_out0,
    output wire [BITNUMBER-1:0] data_out1,
    output wire D0_can_pop,
    output wire D1_can_pop,
	output wire Main_pause
    );


//Wires
wire Main_fifo_full, Main_fifo_empty, Main_Fifo_rd_error, Main_Fifo_wr_error, Main_Fifo_error, Main_almost_full, Main_almost_empty, Main_can_pop,/* Main_pause ,*/ Main_valid_read;
wire VC0_full, VC0_empty, VC0_rd_error, VC0_wr_error, VC0_error, VC0_almost_full, VC0_almost_empty, VC0_can_pop, VC0_pause , VC0_valid_read;
wire VC1_full, VC1_empty, VC1_rd_error, VC1_wr_error, VC1_error, VC1_almost_full, VC1_almost_empty, VC1_can_pop, VC1_pause , VC1_valid_read;
wire D0_full, D0_empty, D0_rd_error, D0_wr_error, D0_error, D0_almost_full, D0_almost_empty, /*D0_can_pop,*/ D0_pause , D0_valid_read;
wire D1_full, D1_empty, D1_rd_error, D1_wr_error, D1_error, D1_almost_full, D1_almost_empty, /*D1_can_pop,*/ D1_pause , D1_valid_read;
wire Mux_valid;
wire pop_main, push_VC0, push_VC1, push_D0, push_D1, pop_VC0, pop_VC1, pop_D0, pop_D1;
wire [BITNUMBER-1:0] Main_Fifo_Data_out, demux_to_VC0, demux_to_VC1, Mux_out, VC0_Data_out, VC1_Data_out, demux_to_D0, demux_to_D1;

fifo #(.BITNUMBER (BITNUMBER), .LENGTH (LENGTH))Main_fifo_(
						      // Outputs
						      .Fifo_full	    (Main_fifo_full),
						      .Fifo_empty	    (Main_fifo_empty),
						      .Fifo_Data_out	(Main_Fifo_Data_out[BITNUMBER-1:0]),
						      .Fifo_rd_error	(Main_Fifo_rd_error),
						      .Fifo_wr_error	(Main_Fifo_wr_error),
						      .Fifo_error	    (Main_Fifo_error),
						      .almost_full	    (Main_almost_full),
						      .almost_empty	    (Main_almost_empty),
						      .can_pop		    (Main_can_pop),
						      .pause		    (Main_pause),
						      .valid_read	    (Main_valid_read),
						      // Inputs
						      .Fifo_Data_in	    (data_in[BITNUMBER-1:0]),
						      .clk		        (clk),
						      .reset		    (reset),
						      .Fifo_rd		    (pop_main),/****/
						      .Fifo_wr		    (push));

demux_id demux_id_(
	// Outputs
    .demux_to_VC0	(demux_to_VC0[BITNUMBER-1:0]),
    .demux_to_VC1	(demux_to_VC1[BITNUMBER-1:0]),
    .Fifo_wr0		(push_VC0),
	.Fifo_wr1		(push_VC1),
	// Inputs
	.Fifo_Data_out 	(Main_Fifo_Data_out[BITNUMBER-1:0]),
    .clk			(clk),
    .reset			(reset),
    .valid_read		(Main_valid_read)
);

fifo #(.BITNUMBER (BITNUMBER), .LENGTH (LENGTH*4))VC0_(
						      // Outputs
						      .Fifo_full	    (VC0_full),
						      .Fifo_empty	    (VC0_empty),
						      .Fifo_Data_out	(VC0_Data_out[BITNUMBER-1:0]),
						      .Fifo_rd_error	(VC0_rd_error),
						      .Fifo_wr_error	(VC0_wr_error),
						      .Fifo_error	    (VC0_error),
						      .almost_full	    (VC0_almost_full),
						      .almost_empty	    (VC0_almost_empty),
						      .can_pop		    (VC0_can_pop),
						      .pause		    (VC0_pause),
						      .valid_read	    (VC0_valid_read),
						      // Inputs
						      .Fifo_Data_in	    (demux_to_VC0[BITNUMBER-1:0]),
						      .clk		        (clk),
						      .reset		    (reset),
						      .Fifo_rd		    (pop_VC0),/****/
						      .Fifo_wr		    (push_VC0));

fifo #(.BITNUMBER (BITNUMBER), .LENGTH (LENGTH*4))VC1_(
						      // Outputs
						      .Fifo_full	    (VC1_full),
						      .Fifo_empty	    (VC1_empty),
						      .Fifo_Data_out	(VC1_Data_out[BITNUMBER-1:0]),
						      .Fifo_rd_error	(VC1_rd_error),
						      .Fifo_wr_error	(VC1_wr_error),
						      .Fifo_error	    (VC1_error),
						      .almost_full	    (VC1_almost_full),
						      .almost_empty	    (VC1_almost_empty),
						      .can_pop		    (VC1_can_pop),
						      .pause		    (VC1_pause),
						      .valid_read	    (VC1_valid_read),
						      // Inputs
						      .Fifo_Data_in	    (demux_to_VC1[BITNUMBER-1:0]),
						      .clk		        (clk),
						      .reset		    (reset),
						      .Fifo_rd		    (pop_VC1),/****/
						      .Fifo_wr		    (push_VC1));

mux_dst #(.BITNUMBER (BITNUMBER))Mux_(
                            // Outputs
                            .valid_out_dest    (Mux_valid),
                            .data_out_dest      (Mux_out[BITNUMBER-1:0]),
                            // Inputs
                            .clk                (clk),
                            .reset              (reset),
                            .data_in0           (VC0_Data_out[BITNUMBER-1:0]),
                            .data_in1           (VC1_Data_out[BITNUMBER-1:0]),
                            .valid_VC0          (VC0_valid_read),
                            .valid_VC1          (VC1_valid_read));

demux_t #(.BITNUMBER (BITNUMBER)) demux_(
                            // Outputs
                            .data_D0        (demux_to_D0[BITNUMBER-1:0]),
                            .data_D1        (demux_to_D1[BITNUMBER-1:0]),
                            .push_D0        (push_D0),
                            .push_D1        (push_D1),
                            // Inputs
                            .clk            (clk), 
                            .reset          (reset),
                            .Mux_out        (Mux_out[BITNUMBER-1:0]),
                            .Mux_valid      (Mux_valid));

fifo #(.BITNUMBER (BITNUMBER), .LENGTH (LENGTH))D0_(
						      // Outputs
						      .Fifo_full	    (D0_full),
						      .Fifo_empty	    (D0_empty),
						      .Fifo_Data_out	(data_out0[BITNUMBER-1:0]),
						      .Fifo_rd_error	(D0_rd_error),
						      .Fifo_wr_error	(D0_wr_error),
						      .Fifo_error	    (D0_error),
						      .almost_full	    (D0_almost_full),
						      .almost_empty	    (D0_almost_empty),
						      .can_pop		    (D0_can_pop),
						      .pause		    (D0_pause),
						      .valid_read	    (D0_valid_read),
						      // Inputs
						      .Fifo_Data_in	    (demux_to_D0[BITNUMBER-1:0]),
						      .clk		        (clk),
						      .reset		    (reset),
						      .Fifo_rd		    (pop_D0),/****/
						      .Fifo_wr		    (push_D0));

fifo #(.BITNUMBER (BITNUMBER), .LENGTH (LENGTH))D1_(
						      // Outputs
						      .Fifo_full	    (D1_full),
						      .Fifo_empty	    (D1_empty),
						      .Fifo_Data_out	(data_out1[BITNUMBER-1:0]),
						      .Fifo_rd_error	(D1_rd_error),
						      .Fifo_wr_error	(D1_wr_error),
						      .Fifo_error	    (D1_error),
						      .almost_full	    (D1_almost_full),
						      .almost_empty	    (D1_almost_empty),
						      .can_pop		    (D1_can_pop),
						      .pause		    (D1_pause),
						      .valid_read	    (D1_valid_read),
						      // Inputs
						      .Fifo_Data_in	    (demux_to_D1[BITNUMBER-1:0]),
						      .clk		        (clk),
						      .reset		    (reset),
						      .Fifo_rd		    (pop_D1),/****/
						      .Fifo_wr		    (push_D1));

assign pop_main = !(VC0_pause || VC1_pause) && !(Main_fifo_empty); // talvez cambiar el !Main_fifo_empty por Main_can_pop
assign pop_VC0 = !(D0_pause || D1_pause) && !(VC0_empty); // VC0_can_pop
assign pop_VC1 = !(D0_pause || D1_pause) && !(VC1_empty); // VC1_can_pop

endmodule
